COL1|COL2
c1|v1
c2|v2